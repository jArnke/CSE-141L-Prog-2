module FourMux #(parameter W=8)(				
	input [1:0] Select,

	input [W-1:0]   A,
			B,
			C,
			D,

	output logic [W-1:0] Out
);


always_comb begin
	Out = A;
	case (Select)
		2'b00: Out = A;
		2'b01: Out = B;
		2'b10: Out = C;
		2'b11: Out = D;
	endcase
end

endmodule